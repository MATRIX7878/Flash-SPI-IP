PACKAGE flashStates IS
    TYPE state IS (INIT, LOADCMD, SEND, LOADADDR, READ, WRITE, DONE);
END PACKAGE;