LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD_UNSIGNED.ALL;

ENTITY conv IS
    PORT(clk : IN STD_LOGIC;
         char : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
         hexLow, hexHigh : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0')
        );
END ENTITY;

ARCHITECTURE behavior OF conv IS
SIGNAL flip : STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');

IMPURE FUNCTION FLIPPER (data : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
VARIABLE var : STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
BEGIN
    FOR i IN 0 TO 7 LOOP
        var(i) := data(7 - i);
    END LOOP;
    RETURN var;
END FUNCTION;

BEGIN
    PROCESS(ALL)
    BEGIN
        IF RISING_EDGE(clk) THEN
            flip <= FLIPPER(char);
            hexLow <= flip(7 DOWNTO 4) + TO_STDLOGICVECTOR(48, 8) WHEN flip(7 DOWNTO 4) <= 9 ELSE flip(7 DOWNTO 4) + TO_STDLOGICVECTOR(55, 8);
            hexHigh <= flip(3 DOWNTO 0) + TO_STDLOGICVECTOR(48, 8) WHEN flip(3 DOWNTO 0) <= 9 ELSE flip(3 DOWNTO 0) + TO_STDLOGICVECTOR(55, 8);
        END IF;
    END PROCESS;
END ARCHITECTURE;
